module scorenumM (
								input [8:0] C_ones,
								input [8:0] C_tens,

								output logic [0:4799] ones,
								output logic [0:4799] tens,
								output logic F_LAG
							 );					 
always_comb 
begin
	F_LAG = 1'b0;
	if(C_ones == 9'b000000000) 
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000111000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000111000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end


	else if((C_ones == 9'b000000001) || (C_ones == 9'b000000010) || (C_ones == 9'b0000000011))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001010000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111100;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if((C_ones == 9'b000000100) || (C_ones == 9'b000000101) || (C_ones == 9'b000000110))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000111000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001001000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111100;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end

	else if((C_ones == 9'b000000111) || (C_ones == 9'b000001000) || (C_ones == 9'b000001001))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011110000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001110000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011111000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end

	else if((C_ones == 9'b000001010) || (C_ones == 9'b000001011) || (C_ones == 9'b000001100))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111100;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end

	else if((C_ones == 9'b000001101) || (C_ones == 9'b000001110) || (C_ones == 9'b000001111))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111100;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000111000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if((C_ones == 9'b000010000) || (C_ones == 9'b000010001) || (C_ones == 9'b000010010))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010111000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011000100;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000100;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end

else if((C_ones == 9'b000010011) || (C_ones == 9'b000010100) || (C_ones == 9'b000010101))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000011111000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end

else if((C_ones == 9'b000010110) || (C_ones == 9'b000010111) || (C_ones == 9'b000011000))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001001000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001001000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000100;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end


else if((C_ones == 9'b000011001) || (C_ones == 9'b000011010) || (C_ones == 9'b000011011))
	begin
	
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001001000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000100;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000001100000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else
	begin
	F_LAG = 1'b1;
	ones[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ones[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	ones[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	ones[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	
	if (C_tens == 9'b000000000)
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000111000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000111000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	else if ((C_tens == 9'b000000001) || (C_tens == 9'b000000010) || (C_tens == 9'b0000000011)) 
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000110000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000001010000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111100000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if ((C_tens == 9'b000000100) || (C_tens == 9'b000000101) || (C_tens == 9'b000000110))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000111000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000001001000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111100000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if ((C_tens == 9'b000000111) || (C_tens == 9'b000001000) || (C_tens == 9'b000001001))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000111100000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000011100000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000111110000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
													
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if ((C_tens == 9'b000001010) || (C_tens == 9'b000001011) || (C_tens == 9'b000001100))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111100000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if ((C_tens == 9'b000001101) || (C_tens == 9'b000001110) || (C_tens == 9'b000001111))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000001111100000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000111000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
		else if ((C_tens == 9'b000010000) || (C_tens == 9'b000010001) || (C_tens == 9'b000010010))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000001111000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000010111000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000011000100000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000010000100000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
		else if ((C_tens == 9'b000010011) || (C_tens == 9'b000010100) || (C_tens == 9'b000010101))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000011111000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if ((C_tens == 9'b000010110) || (C_tens == 9'b000010111) || (C_tens == 9'b000011000))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000110000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000001001000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000110000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000001001000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000010000100000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	else if ((C_tens == 9'b000011001) || (C_tens == 9'b000011010) || (C_tens == 9'b000011011))
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000110000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000001001000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000010000100000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000001111000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000001100000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
	
	
   else
	begin
	
	tens[0:79]       = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[80:159]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[160:239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[240:319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[320:399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[400:479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[480:559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[560:639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[640:719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[720:799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	tens[800:879]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[880:959]      = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[960:1039]     = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1040:1119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1120:1199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1200:1279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1280:1359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1360:1439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1440:1519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1520:1599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[1600:1679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1680:1759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1760:1839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1840:1919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[1920:1999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2000:2079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2080:2159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2160:2239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2240:2319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2320:2399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[2400:2479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2480:2559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2560:2639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2640:2719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2720:2799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2800:2879]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2880:2959]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[2960:3039]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3040:3119]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3120:3199]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[3200:3279]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3280:3359]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3360:3439]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3440:3519]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3520:3599]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3600:3679]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3680:3759]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3760:3839]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3840:3919]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[3920:3999]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	tens[4000:4079]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4080:4159]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4160:4239]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4240:4319]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4320:4399]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4400:4479]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4480:4559]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4560:4639]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4640:4719]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	tens[4720:4799]    = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;

	end
end
endmodule
