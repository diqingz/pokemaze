module my_maps (input [2:0] count,
					  input E_STATE,
					  output logic [3071:0] C_map
					  );


always_comb begin

	if (count == 3'b000)
	begin
	
	C_map[63:0]    = 64'b0;  
	C_map[127:64]   = 64'h0;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]  =64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[383:320] = 64'b0000000000010000001000000000000000000000000000000000000000000000; 
	C_map[447:384] = 64'b0000000000101000010100000000000000000000000000000000000000000000;  
	C_map[511:448] = 64'b0000000001000100100010000000000000000000000000000000000000000000;  
	C_map[575:512] = 64'b0000000010000011000001000000000000000000000000000000000000000000;  
	C_map[639:576] = 64'b0000000100000011000000100000000000000000000000000000000000000000;
	C_map[703:640] = 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[767:704] = 64'b00000;  
	C_map[831:768] = 64'b00000;  
	C_map[895:832] = 64'b00000;  
	C_map[959:896] = 64'b00000;  
	C_map[1023:960] = 64'b00000; 
	C_map[1087:1024] = 64'b00000; 
	C_map[1151:1088] = 64'b00000; 
	C_map[1215:1152] = 64'b00000; 
	C_map[1279:1216] = 64'b00000; 
	C_map[1343:1280] = 64'b00000; 
	C_map[1407:1344] = 64'b00000; 
	C_map[1471:1408] = 64'b00000; 
	C_map[1535:1472] = 64'b00000; 
	C_map[1599:1536] = 64'h00000; 
	C_map[1663:1600] = 64'h00000; 
	C_map[1727:1664] = 64'h00000; 
	C_map[1791:1728] = 64'h00000; 
	C_map[1855:1792] = 64'h00000; 
	C_map[1919:1856] = 64'h00000; 
	C_map[1983:1920] = 64'h00000; 
	C_map[2047:1984] = 64'h00000; 
	C_map[2111:2048] = 64'h00000; 
	C_map[2175:2112] = 64'h00000; 
	C_map[2239:2176] = 64'h00000; 
	C_map[2303:2240] = 64'h00000; 
	C_map[2367:2304] = 64'h00000; 
	C_map[2431:2368] = 64'h00000; 
	C_map[2495:2432] = 64'h00000; 
	C_map[2559:2496] = 64'h00000; 
	C_map[2623:2560] = 64'h00000; 
	C_map[2687:2624] = 64'h00000; 
	C_map[2751:2688] = 64'h00000; 
	C_map[2815:2752] = 64'h00000; 
	C_map[2879:2816] = 64'h00000; 
	C_map[2943:2880] = 64'h00000; 
	C_map[3007:2944] = 64'h00000; 
	C_map[3071:3008] = 64'h00000; 
	
	end
	
	else if (E_STATE)
	begin
	C_map[63:0]    = 64'h00000;  
	C_map[127:64]   = 64'h00000;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]   = 64'b01111011101110100010;  
	C_map[383:320] = 64'b00001010001010110110; 
	C_map[447:384] = 64'b01111001001110101010;  
	C_map[511:448] = 64'b00001000101010100010;  
	C_map[575:512] = 64'b01111011101010100010;  
	C_map[639:576] = 64'h00000;  
	C_map[703:640] = 64'h00000; 
	C_map[767:704] = 64'h00000;  
	C_map[831:768] = 64'h00000;  
	C_map[895:832] = 64'h00000;  
	C_map[959:896] = 64'h00000;  
	C_map[1023:960] = 64'h00000; 
	C_map[1087:1024] = 64'h00000; 
	C_map[1151:1088] = 64'h00000; 
	C_map[1215:1152] = 64'h00000; 
	C_map[1279:1216] = 64'h00000; 
	C_map[1343:1280] = 64'h00000; 
	C_map[1407:1344] = 64'h00000; 
	C_map[1471:1408] = 64'h00000; 
	C_map[1535:1472] = 64'h00000; 
	C_map[1599:1536] = 64'h00000; 
	C_map[1663:1600] = 64'h00000; 
	C_map[1727:1664] = 64'h00000; 
	C_map[1791:1728] = 64'h00000; 
	C_map[1855:1792] = 64'h00000; 
	C_map[1919:1856] = 64'h00000; 
	C_map[1983:1920] = 64'h00000; 
	C_map[2047:1984] = 64'h00000; 
	C_map[2111:2048] = 64'h00000; 
	C_map[2175:2112] = 64'h00000; 
	C_map[2239:2176] = 64'h00000; 
	C_map[2303:2240] = 64'h00000; 
	C_map[2367:2304] = 64'h00000; 
	C_map[2431:2368] = 64'h00000; 
	C_map[2495:2432] = 64'h00000; 
	C_map[2559:2496] = 64'h00000; 
	C_map[2623:2560] = 64'h00000; 
	C_map[2687:2624] = 64'h00000; 
	C_map[2751:2688] = 64'h00000; 
	C_map[2815:2752] = 64'h00000; 
	C_map[2879:2816] = 64'h00000; 
	C_map[2943:2880] = 64'h00000; 
	C_map[3007:2944] = 64'h00000; 
	C_map[3071:3008] = 64'h00000; 
	end
	

	else if (count == 3'b001)
	begin
	C_map[63:0]    = 64'b1111111111111111111111111111111111111111111111111111101110000111;  
	C_map[127:64]  = 64'b0111111111111111111111111110000000000000000000011111111111111111;  
	C_map[191:128] = 64'b1000011100000000000000000000000000000000000000000011111111111111;  
	C_map[255:192] = 64'b1000000000000000000000000000000000000000000000000000000000000111;  
	C_map[319:256] = 64'b0111111111110000000000000000000000000000000000000000000011111111;  
	C_map[383:320] = 64'b1000000000000000000000000000000000000000000000000000000011111111; 
	C_map[447:384] = 64'b0111111111111111111111111111111111111111000000000111111111111111;  
	C_map[511:448] = 64'b1000000000000000000000000000000001111111000000000111111111111111;  
	C_map[575:512] = 64'b1111111111111111111111111111111111111111100000001111111111111111;  
	C_map[639:576] = 64'b0000011111111111111111111111111111100000000000000000000001111111;  
	C_map[703:640] = 64'b1111111111111111111111111111111111100000000000001111111111111111; 
	C_map[767:704] = 64'b1111111111111111111111111111111111100000000000001111111111111111;  
	C_map[831:768] = 64'b1111111111111111111111111111111111100000000000111111111111111111;  
	C_map[895:832] = 64'b1111111111111111111111111111100000000000000000000000001111111111;  
	C_map[959:896] = 64'b1111111111111111111111111111000000000000000000011111111111100000;  
	C_map[1023:960] = 64'b111111111111111111111111111000000000000000000011111111111111111; 
	C_map[1087:1024] = 64'b00000; 
	C_map[1151:1088] = 64'b00000; 
	C_map[1215:1152] = 64'b00000; 
	C_map[1279:1216] = 64'b00000; 
	C_map[1343:1280] = 64'b00000; 
	C_map[1407:1344] = 64'b00000; 
	C_map[1471:1408] = 64'b00000; 
	C_map[1535:1472] = 64'b00000; 
	C_map[1599:1536] = 64'b00000; 
	C_map[1663:1600] = 64'b00000; 
	C_map[1727:1664] = 64'b00000; 
	C_map[1791:1728] = 64'b00000; 
	C_map[1855:1792] = 64'b00000; 
	C_map[1919:1856] = 64'b00000; 
	C_map[1983:1920] = 64'b00000; 
	C_map[2047:1984] = 64'b00000; 
	C_map[2111:2048] = 64'b00000; 
	C_map[2175:2112] = 64'b00000; 
	C_map[2239:2176] = 64'b00000; 
	C_map[2303:2240] = 64'b00000; 
	C_map[2367:2304] = 64'b00000; 
	C_map[2431:2368] = 64'b00000; 
	C_map[2495:2432] = 64'b00000; 
	C_map[2559:2496] = 64'b00000; 
	C_map[2623:2560] = 64'b00000; 
	C_map[2687:2624] = 64'b00000; 
	C_map[2751:2688] = 64'b00000; 
	C_map[2815:2752] = 64'b00000; 
	C_map[2879:2816] = 64'b00000; 
	C_map[2943:2880] = 64'b00000; 
	C_map[3007:2944] = 64'b00000; 
	C_map[3071:3008] = 64'b00000; 
	 
	end
	
	else if (count == 3'b010)
	begin						  
	C_map[63:0]    = 64'h00000;  
	C_map[127:64]   = 64'h00000;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]   = 64'b0;  
	C_map[383:320] = 64'b0000; 
	C_map[447:384] = 64'b00;  
	C_map[511:448] = 64'b00;  
	C_map[575:512] = 64'b00;  
	C_map[639:576] = 64'h00000;  
	C_map[703:640] = 64'h00000; 
	C_map[767:704] = 64'h00000;  
	C_map[831:768] = 64'h00000;  
	C_map[895:832] = 64'h00000;  
	C_map[959:896] = 64'h00000;  
	C_map[1023:960] = 64'h00000; 
	C_map[1087:1024] = 64'h00000; 
	C_map[1151:1088] = 64'h00000; 
	C_map[1215:1152] = 64'h00000; 
	C_map[1279:1216] = 64'h00000; 
	C_map[1343:1280] = 64'h00000; 
	C_map[1407:1344] = 64'h00000; 
	C_map[1471:1408] = 64'h00000; 
	C_map[1535:1472] = 64'h00000; 
	C_map[1599:1536] = 64'h00000; 
	C_map[1663:1600] = 64'h00000; 
	C_map[1727:1664] = 64'h00000; 
	C_map[1791:1728] = 64'h00000; 
	C_map[1855:1792] = 64'h00000; 
	C_map[1919:1856] = 64'h00000; 
	C_map[1983:1920] = 64'h00000; 
	C_map[2047:1984] = 64'h00000; 
	C_map[2111:2048] = 64'h00000; 
	C_map[2175:2112] = 64'h00000; 
	C_map[2239:2176] = 64'h00000; 
	C_map[2303:2240] = 64'h00000; 
	C_map[2367:2304] = 64'h00000; 
	C_map[2431:2368] = 64'h00000; 
	C_map[2495:2432] = 64'h00000; 
	C_map[2559:2496] = 64'h00000; 
	C_map[2623:2560] = 64'h00000; 
	C_map[2687:2624] = 64'h00000; 
	C_map[2751:2688] = 64'h00000; 
	C_map[2815:2752] = 64'h00000; 
	C_map[2879:2816] = 64'h00000; 
	C_map[2943:2880] = 64'h00000; 
	C_map[3007:2944] = 64'h00000; 
	C_map[3071:3008] = 64'h00000;
	end
	
	else if (count == 3'b011)
	begin
	C_map[63:0]    = 64'h00000;  
	C_map[127:64]   = 64'h00000;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]   = 64'b01111011101110100010;  
	C_map[383:320] = 64'b00001010001010110110; 
	C_map[447:384] = 64'b01111001001110101010;  
	C_map[511:448] = 64'b00001000101010100010;  
	C_map[575:512] = 64'b01111011101010100010;  
	C_map[639:576] = 64'h00000;  
	C_map[703:640] = 64'h00000; 
	C_map[767:704] = 64'h00000;  
	C_map[831:768] = 64'h00000;  
	C_map[895:832] = 64'h00000;  
	C_map[959:896] = 64'h00000;  
	C_map[1023:960] = 64'h00000; 
	C_map[1087:1024] = 64'h00000; 
	C_map[1151:1088] = 64'h00000; 
	C_map[1215:1152] = 64'h00000; 
	C_map[1279:1216] = 64'h00000; 
	C_map[1343:1280] = 64'h00000; 
	C_map[1407:1344] = 64'h00000; 
	C_map[1471:1408] = 64'h00000; 
	C_map[1535:1472] = 64'h00000; 
	C_map[1599:1536] = 64'h00000; 
	C_map[1663:1600] = 64'h00000; 
	C_map[1727:1664] = 64'h00000; 
	C_map[1791:1728] = 64'h00000; 
	C_map[1855:1792] = 64'h00000; 
	C_map[1919:1856] = 64'h00000; 
	C_map[1983:1920] = 64'h00000; 
	C_map[2047:1984] = 64'h00000; 
	C_map[2111:2048] = 64'h00000; 
	C_map[2175:2112] = 64'h00000; 
	C_map[2239:2176] = 64'h00000; 
	C_map[2303:2240] = 64'h00000; 
	C_map[2367:2304] = 64'h00000; 
	C_map[2431:2368] = 64'h00000; 
	C_map[2495:2432] = 64'h00000; 
	C_map[2559:2496] = 64'h00000; 
	C_map[2623:2560] = 64'h00000; 
	C_map[2687:2624] = 64'h00000; 
	C_map[2751:2688] = 64'h00000; 
	C_map[2815:2752] = 64'h00000; 
	C_map[2879:2816] = 64'h00000; 
	C_map[2943:2880] = 64'h00000; 
	C_map[3007:2944] = 64'h00000; 
	C_map[3071:3008] = 64'h00000; 
	end
	
	else
	begin
	C_map[63:0]    = 64'h00000;  
	C_map[127:64]   = 64'h00000;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]   = 64'b01111011101110100010;  
	C_map[383:320] = 64'b00001010001010110110; 
	C_map[447:384] = 64'b01111001001110101010;  
	C_map[511:448] = 64'b00001000101010100010;  
	C_map[575:512] = 64'b01111011101010100010;  
	C_map[639:576] = 64'h00000;  
	C_map[703:640] = 64'h00000; 
	C_map[767:704] = 64'h00000;  
	C_map[831:768] = 64'h00000;  
	C_map[895:832] = 64'h00000;  
	C_map[959:896] = 64'h00000;  
	C_map[1023:960] = 64'h00000; 
	C_map[1087:1024] = 64'h00000; 
	C_map[1151:1088] = 64'h00000; 
	C_map[1215:1152] = 64'h00000; 
	C_map[1279:1216] = 64'h00000; 
	C_map[1343:1280] = 64'h00000; 
	C_map[1407:1344] = 64'h00000; 
	C_map[1471:1408] = 64'h00000; 
	C_map[1535:1472] = 64'h00000; 
	C_map[1599:1536] = 64'h00000; 
	C_map[1663:1600] = 64'h00000; 
	C_map[1727:1664] = 64'h00000; 
	C_map[1791:1728] = 64'h00000; 
	C_map[1855:1792] = 64'h00000; 
	C_map[1919:1856] = 64'h00000; 
	C_map[1983:1920] = 64'h00000; 
	C_map[2047:1984] = 64'h00000; 
	C_map[2111:2048] = 64'h00000; 
	C_map[2175:2112] = 64'h00000; 
	C_map[2239:2176] = 64'h00000; 
	C_map[2303:2240] = 64'h00000; 
	C_map[2367:2304] = 64'h00000; 
	C_map[2431:2368] = 64'h00000; 
	C_map[2495:2432] = 64'h00000; 
	C_map[2559:2496] = 64'h00000; 
	C_map[2623:2560] = 64'h00000; 
	C_map[2687:2624] = 64'h00000; 
	C_map[2751:2688] = 64'h00000; 
	C_map[2815:2752] = 64'h00000; 
	C_map[2879:2816] = 64'h00000; 
	C_map[2943:2880] = 64'h00000; 
	C_map[3007:2944] = 64'h00000; 
	C_map[3071:3008] = 64'h00000; 
	end
	
//
//	if (count == 3'b000)
//	begin
//	C_map[19:0]    = 20'h00000;  
//	C_map[39:20]   = 20'h00000;  
//	C_map[59:40]   = 20'h00000;  
//	C_map[79:60]   = 20'h00000;  
//	C_map[99:80]   = 20'b01111011101110100010;  
//	C_map[119:100] = 20'b00001010001010110110; 
//	C_map[139:120] = 20'b01111001001110101010;  
//	C_map[159:140] = 20'b00001000101010100010;  
//	C_map[179:160] = 20'b01111011101010100010;  
//	C_map[199:180] = 20'h00000;  
//	C_map[219:200] = 20'h00000; 
//	C_map[239:220] = 20'h00000;  
//	C_map[259:240] = 20'h00000;  
//	C_map[279:260] = 20'h00000;  
//	C_map[299:280] = 20'h00000;  
//	end
//	
//	else if (E_STATE)
//	begin
//	C_map[19:0]    = 20'h00000;  
//	C_map[39:20]   = 20'h00000;  
//	C_map[59:40]   = 20'h00000;  
//	C_map[79:60]   = 20'h00000;  
//	C_map[99:80]   = 20'h00000;  
//	C_map[119:100] = 20'b00111000100010001110; 
//	C_map[139:120] = 20'b01001000100110000010;  
//	C_map[159:140] = 20'b01001000101010001110;  
//	C_map[179:160] = 20'b01001000110010000010;  
//	C_map[199:180] = 20'b00111000100010001110; 
//	C_map[219:200] = 20'h00000; 
//	C_map[239:220] = 20'h00000;  
//	C_map[259:240] = 20'h00000;  
//	C_map[279:260] = 20'h00000;  
//	C_map[299:280] = 20'h00000;  
//	end
//	
//
//	else if (count == 3'b001)
//	begin
//	C_map[19:0]    = 20'b11111111111111111111;  
//	C_map[39:20]   = 20'b11111110001111111111;  
//	C_map[59:40]   = 20'b00000110000000011000;  
//	C_map[79:60]   = 20'b00000111111100011110;  
//	C_map[99:80]   = 20'b00000111111100011110;  
//	C_map[119:100] = 20'b00000110000000000110;  
//	C_map[139:120] = 20'b00000110011111111110;  
//	C_map[159:140] = 20'b00000110011111111110;  
//	C_map[179:160] = 20'b00000110011000000001; 
//	C_map[199:180] = 20'b00000110000001110001;  
//	C_map[219:200] = 20'b00000111111110000001;  
//	C_map[239:220] = 20'b00000110000000000001;  
//	C_map[259:240] = 20'b11111110011111111111;  
//	C_map[279:260] = 20'b10000000000000000011;  
//	C_map[299:280] = 20'b11111111111111111111;  
//	end
//	
//	else if (count == 3'b010)
//	begin						  
//	C_map[19:0]    = 20'b11111111111111111111;  
//	C_map[39:20]   = 20'b10000000000000000111;  
//	C_map[59:40]   = 20'b11111001110011111111;  
//	C_map[79:60]   = 20'b00001000000011000001;  
//	C_map[99:80]   = 20'b00001001111111011001;  
//	C_map[119:100] = 20'b00001000000011011001;  
//	C_map[139:120] = 20'b00001000111000011001;  
//	C_map[159:140] = 20'b00001111101111111001;  
//	C_map[179:160] = 20'b00000000000000011001;  
//	C_map[199:180] = 20'b11111111111111111001;  
//	C_map[219:200] = 20'b11000000000000000001;  
//	C_map[239:220] = 20'b11101111111111111111;  
//	C_map[259:240] = 20'b11000000000000000011;  
//	C_map[279:260] = 20'b11000000000000000011; 
//	C_map[299:280] = 20'b11111111111111111111; 
//	end
//	
//	else if (count == 3'b011)
//	begin
//	C_map[19:0]    = 20'h00000;  
//	C_map[39:20]   = 20'h00000;  
//	C_map[59:40]   = 20'h0FF00; 
//	C_map[79:60]   = 20'h00900;  
//	C_map[99:80]   = 20'h00900;  
//	C_map[119:100] = 20'h00020;  
//	C_map[139:120] = 20'h00000;  
//	C_map[159:140] = 20'h00000; 
//	C_map[179:160] = 20'h00000;  
//	C_map[199:180] = 20'h00000;  
//	C_map[219:200] = 20'h00000;  
//	C_map[239:220] = 20'h00FF0;  
//	C_map[259:240] = 20'h0F000;  
//	C_map[279:260] = 20'h00000;  
//	C_map[299:280] = 20'h00000; 
//	end
//	
//	else
//	begin
//	C_map[19:0]    = 20'h00000;  
//	C_map[39:20]   = 20'h00000; 
//	C_map[59:40]   = 20'h00000;  
//	C_map[79:60]   = 20'h00000;  
//	C_map[99:80]   = 20'h00000; 
//	C_map[119:100] = 20'b00111000100010001110;  
//	C_map[139:120] = 20'b01001000100110000010;  
//	C_map[159:140] = 20'b01001000101010001110;  
//	C_map[179:160] = 20'b01001000110010000010;  
//	C_map[199:180] = 20'b00111000100010001110;  
//	C_map[219:200] = 20'h00000;  
//	C_map[239:220] = 20'h00000; 
//	C_map[259:240] = 20'h00000;  
//	C_map[279:260] = 20'h00000;  
//	C_map[299:280] = 20'h00000;  
//	end
//	
	
end

endmodule

