module bitmap (input [2:0] count,
					  input E_STATE,
					  input menu_screen,
					  output logic [3071:0] C_map
					  );


always_comb begin

	if (count == 3'b000)
	begin
	
C_map[63:0]    = 64'b0;  
	C_map[127:64]   = 64'h0;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]  = 64'b0000000000000000000000000000000001000000000000000000000000000000;  
	C_map[383:320] =  64'b0000000000000000000000000000000010000000000000000000000000000000; 
	C_map[447:384] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[511:448] =  64'b0000000000000000000000000000000111111101000000100111110001111100;  
	C_map[575:512] =  64'b0000000000000000000000000000000000000100100000101000001010000010;  
	C_map[639:576] =  64'b0000000000000000000000000000000000000100010000101000001010000010;
	C_map[703:640] =  64'b0000000000000000000000000000000000000100001000101000001010000010; 
	C_map[767:704] =  64'b0000000000000000000000000000000000000100000100101000001010000010;  
	C_map[831:768] =  64'b0000000000000000000000000000000000000100000010101000001001111110;  
	C_map[895:832] =  64'b0011110111111100111110001000100111111100000001101000001000000010;  
	C_map[959:896] =  64'b0100010010000001000001010101010000000100000010101000001000000010;  
	C_map[1023:960] = 64'b0100010001000001111111010010010000000100000100101000001000000010; 
	C_map[1087:1024]= 64'b0011110000100001000001010000010000000100001000101000001000000010; 
	C_map[1151:1088]= 64'b0000010000010001000001010000010000000100010000101000001000000010; 
	C_map[1215:1152]= 64'b0000010000001001000001010000010000000100100000101000001000000010; 
	C_map[1279:1216]= 64'b0111110111111101000001010000010111111101000000100111110000000010; 
	C_map[1343:1280]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[1407:1344]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[1471:1408]= 64'b0000000000000000000000000000011100000100100000010101110000000000; 
	C_map[1535:1472]= 64'b0000000000110011100011001111000010000010101110000100001000000000; 
	C_map[1599:1536]= 64'b0000000001001000010100101001000100000001100001010100001000000000; 
	C_map[1663:1600]= 64'b0000000000101000010110101001001000000010100001010100001000000000; 
	C_map[1727:1664]= 64'b0000000001111011100101100111000111000100101110010101110000000000; 
	C_map[1791:1728]= 64'b0000000000000000000000000001000000000000000000000000000000000000; 
	C_map[1855:1792]= 64'b0000000000000000000000000001000000000000000000000000000000000000; 
	C_map[1919:1856]= 64'b0000000000000010000000000000010011100000000001111100000000000000; 
	C_map[1983:1920]= 64'b0000000000000010011010011000010000010000011000010000000000000000; 
	C_map[2047:1984]= 64'b0000000000001111100110100101111100100000100100010000000000000000; 
	C_map[2111:2048]= 64'b0000000000000010000010110100010001000000100100010000000000000000; 
	C_map[2175:2112]= 64'b0000000000000010000010101100010000111000011000010000000000000000; 
	C_map[2239:2176]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2303:2240]= 64'b0000000000000011000000000001100100100000010101110000000000000000; 
	C_map[2367:2304]= 64'b0000000000000000011000001100000010101110000100001000000000000000; 
	C_map[2431:2368]= 64'b0000000000000000010100010100000001100001010100001000000000000000; 
	C_map[2495:2432]= 64'b0000000000000000010010100100000010100001010100001000000000000000; 
	C_map[2559:2496]= 64'b0000000000000000010001000100000100101110010101110000000000000000; 
	C_map[2623:2560]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2687:2624]= 64'b0000000000000000000000000000001100011000000000000011110000000000;
	C_map[2751:2688]= 64'b0000000000000100010011010011001010101001110100110000010000000000; 
	C_map[2815:2752]= 64'b0000000000000100010100110100101001001000001101001001110000000000; 
	C_map[2879:2816]= 64'b0000000000000100010100010010101000001000000101001000010000000000; 
	C_map[2943:2880]= 64'b0000000000000011100100010111001000001000000100110000010000000000; 
	C_map[3007:2944]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[3071:3008]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	end
	
	else if (E_STATE)
	begin
		C_map[63:0]    = 64'b0; 
	C_map[127:64]   = 64'h0;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[383:320] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[447:384] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[511:448] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[575:512] =  64'b0000000000000000000000000000000000000000000000000000000000000000;    
	C_map[639:576] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[703:640] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[767:704] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[831:768] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[895:832] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[959:896] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[1023:960] = 64'b0000000000000000000000000000000000000000000011111110000000000000; 
	C_map[1087:1024]= 64'b0000000000000000000000000000000000000000000000000001000000000000;
	C_map[1151:1088]= 64'b0000000000000000000000000000000000000000000000000001000000000000;
	C_map[1215:1152]= 64'b0000000000000001111110001110111000111111000000000001000000000000;
	C_map[1279:1216]= 64'b0000000000000010000001010001000101000000100111100001000000000000;
	C_map[1343:1280]= 64'b0000000000000001111111010000000101000000100010000001000000000000; 
	C_map[1407:1344]= 64'b0000000000000000000001010000000101100000100010000001000000000000; 
	C_map[1471:1408]= 64'b0000000000000011111110010000000101011111000001111110000000000000;  
	C_map[1535:1472]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[1599:1536]= 64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[1663:1600]= 64'b0000000000000000000000000000000000000000000111111000000000000000; 
	C_map[1727:1664]= 64'b0000000000000000000000000000000000000000001000000100000000000000; 
	C_map[1791:1728]= 64'b0000000000000000000000000000000000000000001000000100000000000000; 
	C_map[1855:1792]= 64'b0000000000000001111101001111110010000000101000000100000000000000; 
	C_map[1919:1856]= 64'b0000000000000000000011010000001001000001001000000100000000000000; 
	C_map[1983:1920]= 64'b0000000000000000000001001111111000100010001000000100000000000000; 
	C_map[2047:1984]= 64'b0000000000000000000001000000001000010100001000000100000000000000; 
	C_map[2111:2048]= 64'b0000000000000000000001011111110000001000000111111000000000000000; 
	C_map[2175:2112]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2239:2176]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2303:2240]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2367:2304]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2431:2368]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2495:2432]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2559:2496]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2623:2560]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2687:2624]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2751:2688]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2815:2752]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2879:2816]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2943:2880]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[3007:2944]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[3071:3008]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	end
	
	else if (menu_screen && count ==3'b001)
	begin
		C_map[63:0]    = 64'hffffffffffffffff;  
	C_map[127:64]   = 64'hffffffffffffffff;  
	C_map[191:128]   = 64'hffffffffffffffff;  
	C_map[255:192]   = 64'hffffffffffffffff;  
	C_map[319:256]   = 64'hffffffffffffffff;  
	C_map[383:320] = 64'hffffffffffffffff; 
	C_map[447:384] = 64'hffffffffffffffff;  
	C_map[511:448] = 64'hffffffffffffffff;  
	C_map[575:512] = 64'hffffffffffffffff;  
	C_map[639:576] = 64'hffffffffffffffff;  
	C_map[703:640] = 64'hffffffffffffffff; 
	C_map[767:704] = 64'hffffffffffffffff;  
	C_map[831:768] = 64'hffffffffffffffff;  
	C_map[895:832] = 64'hffffffffffffffff;  
	C_map[959:896] = 64'hffffffffffffffff;  
	C_map[1023:960] = 64'hffffffffffffffff; 
	C_map[1087:1024] = 64'hffffffffffffffff; 
	C_map[1151:1088] = 64'hffffffffffffffff; 
	C_map[1215:1152] = 64'hffffffffffffffff; 
	C_map[1279:1216] = 64'hffffffffffffffff; 
	C_map[1343:1280] = 64'hffffffffffffffff; 
	C_map[1407:1344] = 64'hffffffffffffffff; 
	C_map[1471:1408] = 64'hffffffffffffffff; 
	C_map[1535:1472] = 64'hffffffffffffffff; 
	C_map[1599:1536] = 64'hffffffffffffffff; 
	C_map[1663:1600] = 64'hffffffffffffffff; 
	C_map[1727:1664] = 64'hffffffffffffffff; 
	C_map[1791:1728] = 64'hffffffffffffffff; 
	C_map[1855:1792] = 64'hffffffffffffffff; 
	C_map[1919:1856] = 64'hffffffffffffffff; 
	C_map[1983:1920] = 64'hffffffffffffffff; 
	C_map[2047:1984] = 64'hffffffffffffffff; 
	C_map[2111:2048] = 64'hffffffffffffffff; 
	C_map[2175:2112] = 64'hffffffffffffffff; 
	C_map[2239:2176] = 64'hffffffffffffffff; 
	C_map[2303:2240] = 64'hffffffffffffffff; 
	C_map[2367:2304] = 64'hffffffffffffffff; 
	C_map[2431:2368] = 64'hffffffffffffffff; 
	C_map[2495:2432] = 64'hffffffffffffffff; 
	C_map[2559:2496] = 64'hffffffffffffffff; 
	C_map[2623:2560] = 64'hffffffffffffffff; 
	C_map[2687:2624] = 64'hffffffffffffffff; 
	C_map[2751:2688] = 64'hffffffffffffffff; 
	C_map[2815:2752] = 64'hffffffffffffffff; 
	C_map[2879:2816] = 64'hffffffffffffffff; 
	C_map[2943:2880] = 64'hffffffffffffffff; 
	C_map[3007:2944] = 64'hffffffffffffffff; 
	C_map[3071:3008] = 64'hffffffffffffffff; 
	end
	
	else if (count == 3'b001 && !menu_screen)
	begin
	C_map[63:0]    = 64'b1111111111111111111111111111111111111111111111111111111111111111;  
	C_map[127:64]  = 64'b1111111111111111111111111110000000000000000000011111111111111111;  
	C_map[191:128] = 64'b1111111111111111000000000000000000000000000000000011111111111111;  
	C_map[255:192] = 64'b1111111111111111000000000000000000000000000000000011111111111111;  
	C_map[319:256] = 64'b1111111111111111000000000000000000000000000000000000000011111111;  
	C_map[383:320] = 64'b1111111111111111000000000000000000000000000000000000000011111111; 
	C_map[447:384] = 64'b1111111111111111111111111111111111111111000000000111111111111111;  
	C_map[511:448] = 64'b1000000000000000000000000000000001111111000000000111111111111111;  
	C_map[575:512] = 64'b1111111111111111111111111111111111111111000000000111111111111111;  
	C_map[639:576] = 64'b1100000000000000000000000000000000000000000000000111111111111111;  
	C_map[703:640] = 64'b1100000000000000000000000000000000000000000000001111111111111111; 
	C_map[767:704] = 64'b1100000000000000000000000000000000000000000000001111111111111111;  
	C_map[831:768] = 64'b1100000000000000000000000000000000000000000000001111111111111111;  
	C_map[895:832] = 64'b1100000011111111111111111111111111111111111111111111111111111111;  
	C_map[959:896] = 64'b1100000011111111111111111111111111111111111111111111111111100000;  
	C_map[1023:960] = 64'b1100000111111111111111111111111111111111111111111111111111100000; 
	C_map[1087:1024] = 64'b1100000000000000000000000000000000000000000000000000000000111111; 
	C_map[1151:1088] = 64'b1100000000000000000000000000000000000000000000000000000000111111; 
	C_map[1215:1152] = 64'b1100000000000000000000000000000000000000000000000000000000111111; 
	C_map[1279:1216] = 64'b1100000000000000000000000000000000000000000000000000000000111111; 
	C_map[1343:1280] = 64'b1111111111111000000111111111111111111111111111111110000000000001; 
	C_map[1407:1344] = 64'b1000000000011000000110000000000000000001111111111110000000000001; 
	C_map[1471:1408] = 64'b1000000000011000000110000000000000000001111111111110000000000001; 
	C_map[1535:1472] = 64'b1111111111111000000111111111111111111111111111111110000000000001; 
	C_map[1599:1536] = 64'b1111000000000000000000000000000000000000000000000000000000000001; 
	C_map[1663:1600] = 64'b1111000000000000000000000000000000000000000000000000000000000001; 
	C_map[1727:1664] = 64'b1111000000000000000000000000000000000000000000000000000000000001; 
	C_map[1791:1728] = 64'b1111000000000000000000000000000000000000000000000000000000000001; 
	C_map[1855:1792] = 64'b1111000000011111111111111111111111111111111111111111111111111111; 
	C_map[1919:1856] = 64'b1111000000011111111111111111111111111111111111111111111111111111; 
	C_map[1983:1920] = 64'b1100000000011111111111111111111111111111111111111111111111111111; 
	C_map[2047:1984] = 64'b1100000000000000000000000000000000000000000000000000000000000001; 
	C_map[2111:2048] = 64'b1100000000000000000000000000000000000000000000000000000000000001; 
	C_map[2175:2112] = 64'b1100000000000000000000000000000000111111111111111111111111111111; 
	C_map[2239:2176] = 64'b1100000000000000000000000000000000111111111111111111111111111111; 
	C_map[2303:2240] = 64'b1111111111111100000000000000000000000000000000000000000000000011; 
	C_map[2367:2304] = 64'b1111111111111100000000000000000000000000000000000000000000000011; 
	C_map[2431:2368] = 64'b1111111111111100000000000000000000000000000000000000000000000011; 
	C_map[2495:2432] = 64'b1111111111111100000000000000000000000000000000000000000000000011; 
	C_map[2559:2496] = 64'b0000011111111100000000000000000000000000000000000000000000000011; 
	C_map[2623:2560] = 64'b0000011111111100000000000000000000000000000000000000000000000011; 
	C_map[2687:2624] = 64'b0000011111111111111111111111111111111111111111111111110000000011; 
	C_map[2751:2688] = 64'b0000011111111111111111111111111111111111111111111111110000000011; 
	C_map[2815:2752] = 64'b1111111111100000000000000000000000000000000000000000000000000011; 
	C_map[2879:2816] = 64'b1111111111100000000000000000000000000000000000000000000000000011; 
	C_map[2943:2880] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	C_map[3007:2944] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	C_map[3071:3008] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	 
	end
	
	else if (count == 3'b010)
	begin						  
	C_map[63:0]    = 64'b1111111111111111111111111111111111111111111111111111111111111111;  
	C_map[127:64]  = 64'b1111111111111111111111111110000000000000000000011111111111111111;  
	C_map[191:128] = 64'b1111111100000000000000000000000000000000000000000011111111111111;  
	C_map[255:192] = 64'b1111111100000000000000000000000000000000000000000000000000000111;  
	C_map[319:256] = 64'b1111111111110000000000000000000000000000000000000000000011111111;  
	C_map[383:320] = 64'b1111111111110000000000000000000000000000000000000000000011111111; 
	C_map[447:384] = 64'b1111111111111111111111111111111111111111000000000111111111111111;  
	C_map[511:448] = 64'b1000000000000000000000000000000001111111000000000111111111111111;  
	C_map[575:512] = 64'b1111111111111111111111111111111111111111100000001111111111111111;  
	C_map[639:576] = 64'b0000011111111111111111111111111111100000000000000000000001111111;  
	C_map[703:640] = 64'b0000011111111111111111111111111111100000000000001111111111111111; 
	C_map[767:704] = 64'b0000011111111111111111111111111111100000000000001111111111111111;  
	C_map[831:768] = 64'b1111111111111111111111111111111111100000000000111111111111111111;  
	C_map[895:832] = 64'b1111111111111111111111111111100000000000000000000000001111111111;  
	C_map[959:896] = 64'b1111111111111111111111111111000000000000000000011111111111100000;  
	C_map[1023:960] = 64'b111111111111111111111111111000000000000000000011111111111100000; 
	C_map[1087:1024] = 64'b1000000000000000000000000111111100000001111111111000000000000000; 
	C_map[1151:1088] = 64'b1000000000000000001111111111111100000000111111111000000000000000; 
	C_map[1215:1152] = 64'b1000000000000000001111111111111100000001111111111111111111111111; 
	C_map[1279:1216] = 64'b1000000000000000001111111111111100000001111111111111111111111111; 
	C_map[1343:1280] = 64'b1000001111100000000000000000000000000001111111111110000000000001; 
	C_map[1407:1344] = 64'b1000000001100000000000000000000000000001111111111110000000000001; 
	C_map[1471:1408] = 64'b1000000001100000000000000000000000000001111111111110000000000001; 
	C_map[1535:1472] = 64'b1000000001111111111111111111111111111111111111111100000000000001; 
	C_map[1599:1536] = 64'b1000000000000000000000000000000000000000000000000000000011000001; 
	C_map[1663:1600] = 64'b1100000000000000000000000000000000000000000000000000000011000001; 
	C_map[1727:1664] = 64'b1110000000000000000000000000000000000000000000000000000011000001; 
	C_map[1791:1728] = 64'b1111000000000000000000000000000000000000000000000000000011000001; 
	C_map[1855:1792] = 64'b1111111111111111111111111111111111111111111111111111111111000001; 
	C_map[1919:1856] = 64'b1100000000000000000000000000000000000000000000000000000000000001; 
	C_map[1983:1920] = 64'b1100000000000000000000000000000000000000000000000000000000000001; 
	C_map[2047:1984] = 64'b1100000000000000000000000000000000000000000000000000000000000001; 
	C_map[2111:2048] = 64'b1100000000000000000000000000000000000000000000000000000000000001; 
	C_map[2175:2112] = 64'b1111111111000000000001111111111111111111111111111111111111111111; 
	C_map[2239:2176] = 64'b1111111111000000000001111111111111111111111111111111111111111111; 
	C_map[2303:2240] = 64'b0000011110000000000000000000000000000000000000000000000000000011; 
	C_map[2367:2304] = 64'b0000011110000000000000000000000000000000000000000000000000000011; 
	C_map[2431:2368] = 64'b0000011111111111100000000000000000000000000000000000000000000011; 
	C_map[2495:2432] = 64'b0000011111111111100000000000000000000000000000000000000000000011; 
	C_map[2559:2496] = 64'b0000011111111111111111111111111111111111000000000000000000000011; 
	C_map[2623:2560] = 64'b0000011111111111111111111111111111111111000000000000000000000011; 
	C_map[2687:2624] = 64'b0000011111111111111111111111111111111111111111111111110000000011; 
	C_map[2751:2688] = 64'b0000011111111111111111111111111111111111111111111111110000000011; 
	C_map[2815:2752] = 64'b1111111111100000000000000000000000000000000000000000000000000011; 
	C_map[2879:2816] = 64'b1111111111100000000000000000000000000000000000000000000000000011; 
	C_map[2943:2880] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	C_map[3007:2944] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	C_map[3071:3008] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	 
	end
	
	else if (count == 3'b011)
	begin
C_map[63:0]    = 64'b1111111111111111111111111111111111111111111111111111111111111111;  
	C_map[127:64]  = 64'b1111111111111111111111111110000000000000000000011111111111111111;  
	C_map[191:128] = 64'b1111111111111111000000000000000000000000000000000011111111111111;  
	C_map[255:192] = 64'b1111111111111111000000000000000000000000000000000011111111111111;  
	C_map[319:256] = 64'b1111111111111111000000000000000000000000000000000000000011111111;  
	C_map[383:320] = 64'b1111111111111111000000000000000000000000000000000000000011111111; 
	C_map[447:384] = 64'b1111111111111111111111111111111111111111000000000111111111111111;  
	C_map[511:448] = 64'b1100000000100000000000000000000001111111000000000111111111111111;  
	C_map[575:512] = 64'b1100000000111111111111111111111111111111000000000111111111111111;  
	C_map[639:576] = 64'b1100000000000000111110000000000000000000000000000111111111111111;  
	C_map[703:640] = 64'b1100000000000000001000000000000000000000000000001111111111111111; 
	C_map[767:704] = 64'b1100000000000000000000000000000000000000000000001111111111111111;  
	C_map[831:768] = 64'b1100000110000000000000000000000000000000000000001111111111111111;  
	C_map[895:832] = 64'b1100000011111110000000111111111111111111111111111111111111111111;  
	C_map[959:896] = 64'b1100000011111111111111111111111111111111111111111111111111100000;  
	C_map[1023:960] = 64'b1100000111111111111111111111111111111111111111111111111111100000; 
	C_map[1087:1024] = 64'b1100000000110000000000011110000000000000000000000000000000111111; 
	C_map[1151:1088] = 64'b1100000000011000000000001111000000000000000000000000000000111111; 
	C_map[1215:1152] = 64'b1100000000001100000000000000000000000000000000000000000000111111; 
	C_map[1279:1216] = 64'b1100000000000000000000000000000000001111100000000000000000111111; 
	C_map[1343:1280] = 64'b1111111100000000000110000000000111111111111111111110000000000001; 
	C_map[1407:1344] = 64'b1111111110000000000111111100000111111111111111111111000000000001; 
	C_map[1471:1408] = 64'b1111111111000000000111111100000111111100000011111110000000000001; 
	C_map[1535:1472] = 64'b1111111111111111111111111111111111111100000011111110000001100001; 
	C_map[1599:1536] = 64'b1111000000000000000000000000000000000000000000000000000000110001; 
	C_map[1663:1600] = 64'b1111000000000000000000000000000000000000000000000000000000011001; 
	C_map[1727:1664] = 64'b1111000000000000000000000000000000000000000000000000000000001101; 
	C_map[1791:1728] = 64'b1111000000011000000000000000000000000000000000000000000000000111; 
	C_map[1855:1792] = 64'b1111000000011111111111111111000011111111111111111111111111111111; 
	C_map[1919:1856] = 64'b1111000000011111111111111111000011111111111111111111111111111111; 
	C_map[1983:1920] = 64'b1111100000011111111111111111111111111111111111111111111111111111; 
	C_map[2047:1984] = 64'b1111100000011111000000000001111110000000000000000000000001100011; 
	C_map[2111:2048] = 64'b1100000000111111000000000001100110000000000000000000000011000011; 
	C_map[2175:2112] = 64'b1100000001111111000000000001100110000000000000000000000110000011; 
	C_map[2239:2176] = 64'b1100000000011111000000000001100110000000000000000000001100000011; 
	C_map[2303:2240] = 64'b1111100000011111000000000001100110000000111110000000011000000011; 
	C_map[2367:2304] = 64'b1111100000000000000000000001100110000000111110000000110000000011; 
	C_map[2431:2368] = 64'b1111100000000000000000000001111110000000111110000000000000000011; 
	C_map[2495:2432] = 64'b1111100000000000000000000000000000000000111110000000000000000011; 
	C_map[2559:2496] = 64'b1111111000000000011111000000000000000000111110000000000000000011; 
	C_map[2623:2560] = 64'b1111111000000000011111000000000000000000111110000110000000000011; 
	C_map[2687:2624] = 64'b1111111111111111111111111111111111111111111111111111000000000011; 
	C_map[2751:2688] = 64'b1111111111111111111111111111111111111111111111111111100000000011; 
	C_map[2815:2752] = 64'b1111111111100000000000000000000000000000000000000000110000000011; 
	C_map[2879:2816] = 64'b1111111111100000000000000000000000000000000000000000010000000011; 
	C_map[2943:2880] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	C_map[3007:2944] = 64'b0000000000000000000000000000000000000000000000000000000000000011; 
	C_map[3071:3008] = 64'b0000000000000000000000000000000000000000000000000000000000000011;
	end
	
	else
	begin
	C_map[63:0]    = 64'b0; 
	C_map[127:64]   = 64'h0;  
	C_map[191:128]   = 64'h00000;  
	C_map[255:192]   = 64'h00000;  
	C_map[319:256]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[383:320] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[447:384] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[511:448] =  64'b0000000000000000000000000000000000000000000000000000000000000000;  
	C_map[575:512] =  64'b0000000000000000000000000000000000000000000000000000000000000000;    
	C_map[639:576] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[703:640] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[767:704] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[831:768] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[895:832] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[959:896] =  64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[1023:960] = 64'b0000000000000000000000000000000000000000000011111110000000000000; 
	C_map[1087:1024]= 64'b0000000000000000000000000000000000000000000000000001000000000000;
	C_map[1151:1088]= 64'b0000000000000000000000000000000000000000000000000001000000000000;
	C_map[1215:1152]= 64'b0000000000000001111110001110111000111111000000000001000000000000;
	C_map[1279:1216]= 64'b0000000000000010000001010001000101000000100111100001000000000000;
	C_map[1343:1280]= 64'b0000000000000001111111010000000101000000100010000001000000000000; 
	C_map[1407:1344]= 64'b0000000000000000000001010000000101100000100010000001000000000000; 
	C_map[1471:1408]= 64'b0000000000000011111110010000000101011111000001111110000000000000;  
	C_map[1535:1472]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[1599:1536]= 64'b0000000000000000000000000000000000000000000000000000000000000000;
	C_map[1663:1600]= 64'b0000000000000000000000000000000000000000000111111000000000000000; 
	C_map[1727:1664]= 64'b0000000000000000000000000000000000000000001000000100000000000000; 
	C_map[1791:1728]= 64'b0000000000000000000000000000000000000000001000000100000000000000; 
	C_map[1855:1792]= 64'b0000000000000001111101001111110010000000101000000100000000000000; 
	C_map[1919:1856]= 64'b0000000000000000000011010000001001000001001000000100000000000000; 
	C_map[1983:1920]= 64'b0000000000000000000001001111111000100010001000000100000000000000; 
	C_map[2047:1984]= 64'b0000000000000000000001000000001000010100001000000100000000000000; 
	C_map[2111:2048]= 64'b0000000000000000000001011111110000001000000111111000000000000000; 
	C_map[2175:2112]= 64'b0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2239:2176]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2303:2240]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2367:2304]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2431:2368]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2495:2432]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2559:2496]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2623:2560]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2687:2624]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2751:2688]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2815:2752]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2879:2816]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[2943:2880]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[3007:2944]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	C_map[3071:3008]= 64'h0000000000000000000000000000000000000000000000000000000000000000; 
	end
	
end

endmodule

